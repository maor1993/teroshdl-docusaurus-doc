module tb_mytb;

mytb dut(
    .rst_n (rst_n),
    .clk (clk),
);


endmodule
