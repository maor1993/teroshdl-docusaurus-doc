//! @title mymodule design
//! @author terosHDL
module myModule #(
    parameter PARAM1 = 1024 //! number of bytes in fifo
)(
    output reg [1023:0] data,
    input clk,
    input rstn
);
    
endmodule