module alwaysmod (
    input clk
);
    
always @(posedge clk ) begin: myproc
    
end
endmodule