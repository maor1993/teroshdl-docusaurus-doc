//! @title mymodule design
//! @author terosHDL
module myModule (
);
    
endmodule